module SPARE_SRAM3KB (/*AUTOARG*/);

endmodule