module BISR(/*AUTOARG*/);






endmodule